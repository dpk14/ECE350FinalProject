module GameLogicController(registers, frame_rt_clk);

    input frame_rt_clk, registers;

    // reads from different registers at frame rate, compares contents

    // TODO: this may be unnecessary, could be handled by processor completely


endmodule