module bitwise_not(out, data_operand);

    input [31:0] data_operand;

    output [31:0] out;

    not not0(out[0], data_operand[0]);
    not not1(out[1], data_operand[1]);
    not not2(out[2], data_operand[2]);
    not not3(out[3], data_operand[3]);
    not not4(out[4], data_operand[4]);
    not not5(out[5], data_operand[5]);
    not not6(out[6], data_operand[6]);
    not not7(out[7], data_operand[7]);
    not not8(out[8], data_operand[8]);
    not not9(out[9], data_operand[9]);
    not not10(out[10], data_operand[10]);
    not not11(out[11], data_operand[11]);
    not not12(out[12], data_operand[12]);
    not not13(out[13], data_operand[13]);
    not not14(out[14], data_operand[14]);
    not not15(out[15], data_operand[15]);
    not not16(out[16], data_operand[16]);
    not not17(out[17], data_operand[17]);
    not not18(out[18], data_operand[18]);
    not not19(out[19], data_operand[19]);
    not not20(out[20], data_operand[20]);
    not not21(out[21], data_operand[21]);
    not not22(out[22], data_operand[22]);
    not not23(out[23], data_operand[23]);
    not not24(out[24], data_operand[24]);
    not not25(out[25], data_operand[25]);
    not not26(out[26], data_operand[26]);
    not not27(out[27], data_operand[27]);
    not not28(out[28], data_operand[28]);
    not not29(out[29], data_operand[29]);
    not not30(out[30], data_operand[30]);
    not not31(out[31], data_operand[31]);

endmodule